* C:\Users\HP\eSim-Workspace\multiplier\multiplier.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/14/21 20:07:01

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  Net-_U3-Pad1_ Net-_U3-Pad2_ Net-_U3-Pad3_ Net-_U3-Pad4_ Net-_U3-Pad5_ Net-_U3-Pad6_ Net-_U3-Pad7_ Net-_U3-Pad8_ multiply		
U6  a0 a1 b0 b1 Net-_U3-Pad1_ Net-_U3-Pad2_ Net-_U3-Pad3_ Net-_U3-Pad4_ adc_bridge_4		
U7  Net-_U3-Pad5_ Net-_U3-Pad6_ Net-_U3-Pad7_ Net-_U3-Pad8_ out1 out2 out3 out4 dac_bridge_4		
R1  out1 GND resistor		
R2  out2 GND resistor		
R3  out3 GND resistor		
R4  out4 GND resistor		
v1  a0 GND pulse		
v2  a1 GND pulse		
v3  b0 GND pulse		
v4  b1 GND pulse		
U5  a0 plot_v1		
U4  a1 plot_v1		
U2  b0 plot_v1		
U1  b1 plot_v1		
U8  out1 plot_v1		
U9  out2 plot_v1		
U10  out3 plot_v1		
U11  out4 plot_v1		

.end
